// spi_system.v

// Generated using ACDS version 15.1 185

`timescale 1 ps / 1 ps
module spi_system (
	 input CLOCK_50,
    input [3:0] KEY,
    output [7:0] LED,
	 input [1:0] SW,
	 
	 output SS_n,
	 output MOSI,
	 input MISO,
	 output SCLK
);

wire [3:0] key_os;
wire [1:0] sw_os;
wire [3:0] delay;
wire main_clk = CLOCK_50;
wire [7:0] data_out;
wire [31:0] count;

oneshot os (
    .clk (main_clk),
    .edge_sig (KEY),
    .level_sig (key_os)
);

oneshot os2 (
    .clk (main_clk),
    .edge_sig (SW),
    .level_sig (sw_os)
);

delay_ctrl dc (
    .clk (main_clk),
    .faster (key_os[1]),
    .slower (key_os[0]),
    .delay (delay),
    .reset (key_os[3])
);

blinker b (
    .clk (main_clk),
    .delay (delay),
    .led (LED[3:0]),
    .reset (key_os[3]),
    .pause (key_os[2])
);

counter c(
	.clock(main_clk),
	.count(count)
);

assign LED[7:4] = count[29:26];

spi_master spi (
	.sclk_i(main_clk),
	.pclk_i(main_clk),
	.rst_i(KEY[3]),
	.spi_ssel_o(SS_n),
   .spi_sck_o(SCLK),
   .spi_mosi_o(MOSI),
   .spi_miso_i(MISO),
//	.di_req_o(LED[7]),
	.di_i(delay),
	.wren_i(SW[0]),
//	.wr_ack_o(LED[6]),
//	.do_valid_o(LED[5]),
	.do_o(data_out)
);

endmodule
