
module powerlink (
	);	

endmodule
