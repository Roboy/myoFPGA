// pid_controller.v

// Generated using ACDS version 16.1 203

`timescale 1 ps / 1 ps
module pid_controller (
	);

	pid_controller_pid_controller_0 pid_controller_0 (
	);

endmodule
