	component powerlink is
	end component powerlink;

	u0 : component powerlink
		port map (
		);

